{%- block instantiate_deta_lut %}
    calc_deta_lut_{{ obj1|lower }}_{{ obj2|lower }}_bx_{{ bx1 }}_bx_{{ bx2 }}_i: entity work.deta_lut
        generic map(
            N_{{ obj1|upper }}_OBJECTS, N_{{ obj2|upper }}_OBJECTS, ({{ obj1|lower }}_t,{{ obj2|lower }}_t)
        )
        port map(
            deta_calc_{{ obj1|lower }}_{{ obj2|lower }}(bx({{ bx1 }}),bx({{ bx2 }})),
            deta_{{ obj1|lower }}_{{ obj2|lower }}(bx({{ bx1 }}),bx({{ bx2 }}))
        );
{%- endblock instantiate_deta_lut %}
