{%- block instantiate_comparators_muon_charge_corr %}
  {%- set o1 = condition.objects[0] %}
  {%- set o2 = condition.objects[1] %}
    comp_muon_charge_corr_{{ condition.chargeCorrelationMode }}_{{ index }}_i: entity work.comparators_muon_charge_corr
        generic map(
            {{ condition.chargeCorrelationMode }}, CC_{{ condition.chargeCorrelation|upper }}
        )
        port map(
            lhc_clk, 
            cc_{{ condition.chargeCorrelationMode }} => cc_{{ condition.chargeCorrelationMode }}(bx({{ o1.object_handle.bx_offset }}),bx({{ o2.object_handle.bx_offset }})), 
            comp_o_{{ condition.chargeCorrelationMode }} => cc_{{ condition.chargeCorrelationMode }}_{{ index }}
        );
{% endblock instantiate_comparators_muon_charge_corr %}
{# eof #}
